module SUM (S,A,B,Cin);
output S;
input A,B,Cin;
assign S=A^B^Cin;
endmodule

