
module sum(S, A, B);
	output S;
	input A, B;
	xor x1(S, A, B);
endmodule
